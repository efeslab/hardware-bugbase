module ila_0 (
    input logic clk,
    input logic [4095:0] probe0,
    input logic [4095:0] probe1
);

endmodule
